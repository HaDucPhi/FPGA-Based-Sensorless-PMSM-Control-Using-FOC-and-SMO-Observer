--
LIBRARY IEEE; -- THU VIEN CHUAN IEEE
USE IEEE.STD_LOGIC_1164.ALL; -- SU DUNG GOI THU VIEN HO TRO CAC PHEP TOAN LOGIC
USE IEEE.STD_LOGIC_ARITH.ALL; -- SU DUNG GOI THU VIEN HO TRO CAC PHEP TOAN SO HOC TREN KIEU DU LIEU STD_LOGIC_VECTOR
USE IEEE.STD_LOGIC_SIGNED.ALL; -- SU DUNG GOI THU VIEN MO RONG KHA NANG SU LY CAC SO NGUYEN CO DAU KIEU STD_LOGIC_VECTOR
--
LIBRARY LPM; -- THU VIEN KHOI TAO LPM
USE LPM.LPM_COMPONENTS.ALL; -- SU DUNG TAT CA CAC GOI THANH PHAN TRONG THU VIEN LPM

ENTITY PLL IS
PORT(
	CLK,CLK_80N		: IN  STD_LOGIC:='0';
	E_ALPHA,E_BETA		: IN  STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
	THETA			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
	SPEED			: BUFFER STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0')
);
END PLL;

ARCHITECTURE PLL_ARCH OF PLL IS
SIGNAL H_ALPHA,H_BETA	: STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
SIGNAL OM		: STD_LOGIC_VECTOR(31 DOWNTO 0):=X"00007CD6";
SIGNAL E,E1,W,WI	: STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
SIGNAL TETA_TEMP	: STD_LOGIC_VECTOR(31 DOWNTO 0):=X"0001921F";
SIGNAL TT,TP		: STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
SIGNAL ERS		: STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
SIGNAL SD1,SD		: STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
SIGNAL SPEED1		: STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
SIGNAL PI		: STD_LOGIC_VECTOR(31 DOWNTO 0):=X"0001921F";
SIGNAL TS		: STD_LOGIC_VECTOR(31 DOWNTO 0):=X"00000034";
SIGNAL KP		: STD_LOGIC_VECTOR(31 DOWNTO 0):=X"00C80000";
SIGNAL KI		: STD_LOGIC_VECTOR(31 DOWNTO 0):=X"00010000";
--
SIGNAL ADDA, ADDB, ADDRS, MULA, MULB,ADDRB 	 : STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
SIGNAL MULR 					 : STD_LOGIC_VECTOR(63 DOWNTO 0):=(OTHERS => '0');
SIGNAL OVERFLOW,COUT				 : STD_LOGIC;
--
SIGNAL ANGLE				 	 : STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
SIGNAL SIN_T,COS_T			 	 : STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS => '0');
--
    COMPONENT SIN_COS
	PORT(
	CLK			: IN STD_LOGIC := '0';  
	THETA			: IN STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
	SIN_OUT			: OUT STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
	COS_OUT			: OUT STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0')
        );
	END COMPONENT;
BEGIN
U: SIN_COS
PORT MAP(
	CLK => CLK,
	THETA => ANGLE,
	SIN_OUT => SIN_T,
	COS_OUT => COS_T
);
    MULL: LPM_MULT
    GENERIC MAP (
        LPM_WIDTHA         => 32,
        LPM_WIDTHB         => 32,
        LPM_WIDTHP         => 64,
        LPM_REPRESENTATION => "SIGNED",
        LPM_PIPELINE       => 1
    )
    PORT MAP (
        DATAA  => MULA, 
        DATAB  => MULB,
        CLOCK  => CLK,
        RESULT => MULR
    );

    ADDER: LPM_ADD_SUB
    GENERIC MAP(
        LPM_WIDTH          => 32,
        LPM_REPRESENTATION => "SIGNED",
        LPM_PIPELINE       => 1
    )
    PORT MAP(
        DATAA 		=> ADDA,
        DATAB 		=> ADDB,
        CLOCK 		=> CLK,
        RESULT 		=> ADDRB,
	OVERFLOW 	=> OVERFLOW,
	COUT 		=> COUT
    );
PROCESS(CLK,ADDRB)
BEGIN
	IF CLK'EVENT AND CLK = '1' THEN -- XU LY TRAN BO CONG
		IF OVERFLOW = '1' THEN
			IF COUT = '1' THEN
				ADDRS <= X"80000000";
			ELSE
				ADDRS <= X"7FFFFFFF";
			END IF;
		ELSE
			ADDRS <= ADDRB;
		END IF;
	END IF;
END PROCESS;

PLL : BLOCK
SIGNAL CNT   : STD_LOGIC_VECTOR(15 DOWNTO 0):=(OTHERS => '0');
BEGIN
  PROCESS(CLK_80N)
  BEGIN
    IF CLK_80N'EVENT AND CLK_80N = '1' THEN
      CNT <= CNT + X"0001";
      IF CNT = X"0000" THEN             	
        ADDA <= -E_ALPHA;
        ADDB <= H_ALPHA;
      ELSIF CNT = X"0001" THEN
	MULA <= ADDRS;
	MULB <= OM;
      ELSIF CNT = X"0002" THEN
	ADDA <= MULR(46 DOWNTO 15);
	ADDB <= E_ALPHA;
      ELSIF CNT = X"0003" THEN
	H_ALPHA <= ADDRS;	-- H_ALPHA(k+1) = Omega*(H_alpha - E_alpha) + E_alpha
      ELSIF CNT = X"0004" THEN
	ADDA <= H_BETA;
	ADDB <= -E_BETA;
      ELSIF CNT = X"0005" THEN
	MULA <= ADDRS;
	MULB <= OM;
      ELSIF CNT = X"0006" THEN
	ADDA <= MULR(46 DOWNTO 15);
	ADDB <= E_BETA;
      ELSIF CNT = X"0007" THEN
	H_BETA <= ADDRS;	-- H_BETA(k+1) = Omega*(H_BETA - E_ALPHA) + E_BETA
      ELSIF CNT = X"0008" THEN
	ANGLE  <= TETA_TEMP;
      ELSIF CNT = X"0009" THEN
	MULA <= COS_T;
	MULB <= -H_ALPHA;
      ELSIF CNT = X"000A" THEN
	ADDA <= MULR(56 DOWNTO 25);
	MULA <= SIN_T;
	MULB <= -H_BETA;
      ELSIF CNT = X"000B" THEN
	ADDB <= MULR(56 DOWNTO 25);
      ELSIF CNT = X"000C" THEN
	E <= ADDRS;		-- E = -H_ALPHA*COS(THETA) - H_BETA*SIN(THETA)
      ELSIF CNT = X"000D" THEN
	ADDA <= WI;
	MULA <= KI;-- 31Q15
	MULB <= E1; -- 31Q20
      ELSIF CNT = X"000E" THEN
	ADDB <= MULR(51 DOWNTO 20);
      ELSIF CNT = X"000F" THEN
	WI <= ADDRS;
	MULA <= KP; -- 31Q15
	MULB <= E;  -- 31Q20
      ELSIF CNT = X"0010" THEN
	ADDA <= MULR(51 DOWNTO 20);
	ADDB <= WI;
      ELSIF CNT = X"0011" THEN
	W    <= ADDRS;		-- W(k) = KP*E(k) + Ki*E(k-1) + WI(k-1)
      ELSIF CNT = X"0012" THEN
	ADDA <= TETA_TEMP;
	MULA <= TS; -- 31Q20
	MULB <= W;  -- 31Q15
      ELSIF CNT = X"0013" THEN
	ADDB <= MULR(51 DOWNTO 20);
      ELSIF CNT = X"0014" THEN
	TETA_TEMP <= ADDRS;	-- TETA_TEMP(k) = TETA_TEMP(k-1) + Ts*W(k)
	ADDA <= TETA_TEMP;
	ADDB <= PI;
      ELSIF CNT = X"0015" THEN
	TT <= ADDRS;
      ELSIF CNT = X"0016" THEN
	IF TT > X"0003243E" THEN
		TT <= X"00000000";
		TETA_TEMP <= X"FFFE6DE1";
	ELSIF TT < X"00000000" THEN
		TT <= X"00000000";
		TETA_TEMP <= X"0001921F";	
	END IF;
      ELSIF CNT = X"0017" THEN           	
        ADDA <= TT;
        ADDB <= -TP;
      ELSIF CNT = X"0018" THEN
	ERS <= ADDRS;
      ELSIF CNT = X"0019" THEN	
	IF ERS > X"00000CCC" OR ERS < X"FFFFF334" THEN
		SD <= SD1;
	ELSE
		MULA <= ERS;
		MULB <= X"09C40000";
	END IF;
      ELSIF CNT = X"001A" THEN	
	IF ERS > X"00000CCC" OR ERS < X"FFFFF334" THEN
		SD <= SD1;
	ELSE
		SD <= MULR(46 DOWNTO 15);
	END IF;	
      ELSIF CNT = X"001B" THEN             	
        ADDA <= -SD1;
        ADDB <= SPEED;
      ELSIF CNT = X"001C" THEN
	MULA <= ADDRS;
	MULB <= OM;
      ELSIF CNT = X"001D" THEN
	ADDA <= MULR(46 DOWNTO 15);
	ADDB <= SD1;
      ELSIF CNT = X"001E" THEN
	SPEED <= ADDRS;	-- SPEED(k+1) = Omega*(SPEED(k) - SD1) + SD1
      ELSIF CNT = X"0270" THEN
	CNT <= X"0000";
	TP <= TT;
	SD1 <= SD;
	THETA <= TT;	
	E1 <= E;
	END IF;
    END IF;
  END PROCESS;
END BLOCK;

END PLL_ARCH;
